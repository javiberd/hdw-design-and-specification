---------------------------------------------------------------------
--
--  Fichero:
--    lab10.vhd  26/10/2017
--
--    (c) J.M. Mendias
--    Dise�o Autom�tico de Sistemas
--    Facultad de Inform�tica. Universidad Complutense de Madrid
--
--  Prop�sito:
--    Laboratorio 10
--
--  Notas de dise�o:
--
---------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity lab10 is
  port
  (
    rstPb_n  : in std_logic;
    osc      : in std_logic;
    switches : inout std_logic_vector(7 downto 0);
    leds     : inout std_logic_vector(7 downto 0);
    upSegs   : inout std_logic_vector(7 downto 0)
  );
end lab10;

---------------------------------------------------------------------

library unisim;
use unisim.vcomponents.all;
use work.common.all;

architecture syn of lab10 is

  signal clk, rst_n : std_logic;
 
  signal apBus : std_logic_vector(9 downto 0);
  signal dpBus : std_logic_vector(17 downto 0);
  signal inPort, outPort : std_logic_vector(7 downto 0);
  signal interrupt, interrupt_ack : std_logic;
 
  signal wrCE, rdCE : std_logic;
  signal aBus, dBus : std_logic_vector(7 downto 0);
 
  signal wrE1, rdE1, int1 : std_logic;
  signal regSel1 : std_logic_vector(0 downto 0);
  signal dataIn1, dataOut1 : std_logic_vector(7 downto 0);

  signal wrE2, rdE2 : std_logic;
  signal regSel2 : std_logic_vector(0 downto 0);
  signal dataIn2, dataOut2 : std_logic_vector(7 downto 0);

  signal wrE3, rdE3 : std_logic;
  signal regSel3 : std_logic_vector(0 downto 0);
  signal dataIn3, dataOut3 : std_logic_vector(7 downto 0);
  
begin

  clk <= osc;
  
  resetSyncronizer : synchronizer
    generic map ( STAGES => 2, INIT => '0' )
    port map ( rst_n => rstPb_n, clk => clk, x => '1', xSync => rst_n );

  ------------------  
 
  gpioWrapper1 : busWrapper
    generic map ( NUMREG => 2, DWIDTH => 8, AWIDTH => 8, BASEADDR => 16#fe# )
    port map ( 
      wrCE => wrCE, rdCE => rdCE, aBus => aBus, dBus => dBus, 
      regSel => regSel1, wrE => wrE1, dataIn => dataIn1, rdE => rdE1, dataOut => dataOut1 
    );

  gpio1 : gpio
    generic map ( DWIDTH => 8, PWIDTH => 8 )
    port map ( 
      rst_n => rst_n, clk => clk, 
      regSel => regSel1(0), wrE => wrE1, dataIn => dataIn1, rdE => rdE1, dataOut => dataOut1, int => int1,
      io => switches 
    ); 

  gpioWrapper2 : busWrapper
    generic map ( NUMREG => 2, DWIDTH => 8, AWIDTH => 8, BASEADDR => 16#fc# )
    port map ( 
      wrCE => wrCE, rdCE => rdCE, aBus => aBus, dBus => dBus, 
      regSel => regSel2, wrE => wrE2, dataIn => dataIn2, rdE => rdE2, dataOut => dataOut2
    );
    
  gpio2 : gpio
    generic map ( DWIDTH => 8, PWIDTH => 8 )
    port map ( 
      rst_n => rst_n, clk => clk, 
      regSel => regSel2(0), wrE => wrE2, dataIn => dataIn2, rdE => rdE2, dataOut => dataOut2, int => open, 
      io => leds
    );

  gpioWrapper3 : busWrapper
    generic map ( NUMREG => 2, DWIDTH => 8, AWIDTH => 8, BASEADDR => 16#fa# )
    port map ( 
      wrCE => wrCE, rdCE => rdCE, aBus => aBus, dBus => dBus, 
      regSel => regSel3, wrE => wrE3, dataIn => dataIn3, rdE => rdE3, dataOut => dataOut3
    );
    
  gpio3 : gpio
    generic map ( DWIDTH => 8, PWIDTH => 8 )
    port map ( 
      rst_n => rst_n, clk => clk, 
      regSel => regSel3(0), wrE => wrE3, dataIn => dataIn3, rdE => rdE3, dataOut => dataOut3, int => open, 
      io => upSegs
    );
     
  intFF:
  process (rst_n, clk)
  begin
    if rst_n='0' then
      interrupt <= '0';
    elsif rising_edge(clk) then
      if int1='1' then
        interrupt <= '1';
      elsif interrupt_ack='1' then
        interrupt <= '0';
      end if;
    end if;
  end process;
  
  microcontroller: kcpsm3
    port map( 
      reset => not rst_n, clk => clk,
      interrupt => interrupt, interrupt_ack => interrupt_ack,
      address => apBus, 
      instruction => dpBus, 
      port_id => aBus, 
      write_strobe => wrCE, out_port => outPort, 
      read_strobe => rdCE, in_port => dBus  
    );   
    
  dBus <= outPort when wrCE='1' else (others => 'Z');
 
  -- Esta memoria contiene el programa memlab10.psm compilado, el cual:
  --   Indefinidamente muestra los numeros 0-f en el display 7-segs conectado al GPIO-3
  --   Cada vez que el procesador recibe una interrupci�n (por un cambio de estado de los switches), escribe en los leds (conectados al GPIO-2) el valor leido en los switches (conectados al GPIO-1)
  programMemory : RAMB16_S18
    generic map (
      INIT_00 => X"01FF80016F3FCFFC4FFEEF3F4005A00F8001000F00430000C00100200019C000",
      INIT_01 => X"A000CFFB0F00CFFD0F00CFFF0FFFA0005410C1015411C2015412C30103FF02FF",
      INIT_02 => X"EF060F5FEF050F5BEF040F33EF030F79EF020F6DEF010F30EF000F7ECFFA0F00",
      INIT_03 => X"EF0E0F4FEF0D0F3DEF0C0F4EEF0B0F1FEF0A0F77EF090F7BEF080F7FEF070F70",
      INIT_04 => X"0000000000000000000000000000000000000000A000CFFA7F00A000EF0F0F47",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"400A000000000000000000000000000000000000000000000000000000000000",
      INITP_00 => X"00000000000000000000000000000A288888888888888888A222DDD0322C7CFF",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"C000000000000000000000000000000000000000000000000000000000000000"
    )  
    port map (
      clk => clk, en => '1', ssr => '0', we => '0',
      addr => apBus,
      di => X"0000", dip => "00",
      do => dpBus(15 downto 0), dop => dpBus(17 downto 16)   
    );
            
end syn;
